module sudoku_v(enter,out,done);
	input [80:0] enter;
	output [80:0] out;
	output done;
	
	
	
endmodule 